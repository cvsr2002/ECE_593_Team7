package riscv_test_pkg;

  import opcodes::*;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "exec_record.svh"
  `include "iss_class.svh"
  `include "execute_driver.svh"
  `include "riscv_monitor.svh"
  `include "execute_agent.svh"
  `include "cpu_tracer.svh"
  `include "execute_scoreboard.svh"
  `include "env_execute_test.svh"
  `include "execute_test.svh"
  `include "mem_test.svh"
  `include "fibonacci.svh"
  
endpackage
