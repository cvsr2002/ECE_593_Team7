
package riscv_opcode_test_pkg;

  import opcodes::*;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "exec_record.svh"
  `include "iss_class.svh"
  `include "riscv_monitor.svh"
  `include "cpu_tracer.svh"
  `include "execute_scoreboard.svh"
  `include "opcode_seq_item.svh"
  `include "opcode_seq.svh"
  `include "opcode_sequencer.svh"
  `include "opcode_driver.svh"
  `include "opcode_agent.svh"
  `include "opcode_env.svh"
  `include "opcode_test.svh"
  
endpackage
